`timescale 1ns / 1ps

module Cell(
    input clk,
    input Sel,
    input Turn,
    input Reset,
    output reg [1:0] State
);

    // Define state encoding
    localparam N = 2'b00, X = 2'b01, O = 2'b11;

    reg [1:0] PS, NS;

    // State register
    always @(posedge clk or posedge Reset) begin
        if (Reset)
            PS <= N;
        else
            PS <= NS;
    end

    // Next-state logic
    always @(*) begin
        case (PS)
            N: begin
                State = 2'b00;
                if (Sel && ~Turn)
                    NS = X;
                else if (Sel && Turn)
                    NS = O;
                else
                    NS = PS;
            end
            X: begin
                State = 2'b01;
                NS = PS;
            end
            O: begin
                State = 2'b11;
                NS = PS;
            end
            default: begin
                State = 2'b00;
                NS = N;
            end
        endcase
    end

endmodule

